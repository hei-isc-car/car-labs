ARCHITECTURE sim OF xor2 IS
BEGIN
  xorOut <= in1 xor in2 after delay;
END ARCHITECTURE sim;
