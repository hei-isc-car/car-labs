ARCHITECTURE sim OF transSignedUlog IS
BEGIN
  out1 <= std_ulogic_vector(in1) after delay;
END ARCHITECTURE sim;
