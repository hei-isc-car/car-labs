ARCHITECTURE sim OF and3 IS
BEGIN
  out1 <= in1 and in2 and in3 after delay;
END ARCHITECTURE sim;
