ARCHITECTURE sim OF onesUnsigned IS
BEGIN
  ones <= (others => '1');
END sim;
