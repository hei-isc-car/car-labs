ARCHITECTURE sim OF onesSigned IS
BEGIN
  ones <= (others => '1');
END sim;
