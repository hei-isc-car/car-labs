ARCHITECTURE sim OF xor5 IS
BEGIN
  xorOut <= in1 xor in2 xor in3 xor in4 xor in5 after delay;
END ARCHITECTURE sim;
