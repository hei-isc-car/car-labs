ARCHITECTURE sim OF logic1 IS
BEGIN
  logic_1 <= '1';
END sim;
