ARCHITECTURE sim OF or5_m IS
BEGIN
  out1 <= in1 or in2 or in3 or in4 or in5 after delay;
END ARCHITECTURE sim;
