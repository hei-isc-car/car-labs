ARCHITECTURE sim OF bufferUnsigned IS
BEGIN
  out1 <= in1 after delay;
END ARCHITECTURE sim;
