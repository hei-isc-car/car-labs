ARCHITECTURE sim OF or2 IS
BEGIN
  out1 <= in1 or in2 after delay;
END ARCHITECTURE sim;
