ARCHITECTURE sim OF or2_m IS
BEGIN
  out1 <= in1 or in2 after delay;
END ARCHITECTURE sim;
