ARCHITECTURE sim OF logic0 IS
BEGIN
  logic_0 <= '0';
END sim;
