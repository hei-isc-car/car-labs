ARCHITECTURE sim OF and2 IS
BEGIN
  out1 <= in1 and in2 after delay;
END ARCHITECTURE sim;
