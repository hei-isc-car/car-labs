ARCHITECTURE sim OF bufferUlogicVector IS
BEGIN
  out1 <= in1 after delay;
END ARCHITECTURE sim;
