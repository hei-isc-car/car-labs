ARCHITECTURE sim OF bufferUlogic IS
BEGIN
  out1 <= in1 after delay;
END ARCHITECTURE sim;
