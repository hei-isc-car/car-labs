LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE gates IS

--  constant gateDelay: time := 1 ns;
  constant gateDelay: time := 0.1 ns;

END gates;
