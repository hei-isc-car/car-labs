ARCHITECTURE sim OF zeroSigned IS
BEGIN
  zero <= (others => '0');
END sim;
