ARCHITECTURE sim OF and4 IS
BEGIN
  out1 <= in1 and in2 and in3 and in4 after delay;
END ARCHITECTURE sim;
