ARCHITECTURE sim OF or4_m IS
BEGIN
  out1 <= in1 or in2 or in3 or in4 after delay;
END ARCHITECTURE sim;
