ARCHITECTURE sim OF xor3 IS
BEGIN
  xorOut <= in1 xor in2 xor in3 after delay;
END ARCHITECTURE sim;
