ARCHITECTURE sim OF subUnsigned IS
BEGIN
  out1 <= in1 - in2 after delay;
END ARCHITECTURE sim;
