ARCHITECTURE sim OF xor4 IS
BEGIN
  xorOut <= in1 xor in2 xor in3 xor in4 after delay;
END ARCHITECTURE sim;
