FILE_NAMING_RULE: %(entity_name)_entity.vhd
DESCRIPTION_START
This is the default template used for the creation of VHDL Entity files.
Template supplied by Mentor Graphics.
DESCRIPTION_END
--
-- VHDL Entity %(library).%(unit).%(view)
--
-- Created:
--          by - %(user).%(group) (%(host))
--          at - %(time) %(date)
--
-- using Mentor Graphics HDL Designer(TM) %(version)
--
%(entity)
