ARCHITECTURE sim OF or3 IS
BEGIN
  out1 <= in1 or in2 or in3 after delay;
END ARCHITECTURE sim;
