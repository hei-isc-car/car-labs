ARCHITECTURE sim OF transLogUlog IS
BEGIN
  out1 <= std_ulogic_vector(in1) after delay;
END ARCHITECTURE sim;
