ARCHITECTURE sim OF and5 IS
BEGIN
  out1 <= in1 and in2 and in3 and in4 and in5 after delay;
END ARCHITECTURE sim;
