FILE_NAMING_RULE: %(entity_name)_%(arch_name).vhd
DESCRIPTION_START
This is the default template used for the creation of combined VHDL Architecture and Entity files.
Template supplied by Mentor Graphics.
DESCRIPTION_END
--
-- VHDL Architecture %(library).%(unit).%(view)
--
-- Created:
--          by - %(user).%(group) (%(host))
--          at - %(time) %(date)
--
-- using Mentor Graphics HDL Designer(TM) %(version)
--
%(entity)
--
%(architecture)
