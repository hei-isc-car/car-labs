ARCHITECTURE sim OF transUnsignedSigned IS
BEGIN
  out1 <= signed(in1) after delay;
END ARCHITECTURE sim;
