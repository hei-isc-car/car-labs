ARCHITECTURE sim OF transSignedUnsigned IS
BEGIN
  out1 <= unsigned(in1) after delay;
END ARCHITECTURE sim;
