ARCHITECTURE sim OF zeroUnsigned IS
BEGIN
  zero <= (others => '0');
END sim;
